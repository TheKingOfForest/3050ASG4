
`timescale 100fs/100fs
module cpu_test;


endmodule